`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/04/11 16:17:19
// Design Name: 
// Module Name: Mult
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Mult#(
    parameter BITWIDTH = 32
)(
    input [BITWIDTH - 1:0] a,
    input [BITWIDTH - 1:0] b,
    input clk,
    output [BITWIDTH - 1:0] c
);
    FLOAT32_MUL_PIPELINE chip (
        .a(a), .b(b), .out(c),
        .clk(clk)
    );
endmodule
