module conv1_params (
    output [32 * 2 * 2 * 3 * 8 - 1 : 0] weight,
    output [32 * 8 - 1 : 0] bias
);
    assign weight = {32'b0111111000011100111001010011101,32'b1111110100100010100011011111101,32'b0111111010000110001001110100101,32'b0111111000011011010010111011001,32'b0111110100111110010111110010010,32'b0111111001000110110110101011000,32'b0111110000001011010000101111111,32'b1111110001110110101000001001110,32'b0111110100001101011111001101011,32'b0111111001011100101010001111100,32'b0111110101001111101110110111000,32'b1111111000101011001111010111110,32'b1111110110110011011101110101010,32'b0111111000011000011111101111100,32'b0111111001011000011010110011101,32'b0111111010011001110110101001111,32'b0111111000111010111010101011011,32'b0111111001101000101101010101111,32'b0111110111110001110000001100100,32'b1111110000100111000011001100111,32'b1111111011000110100100010111100,32'b0111111011000001010110011110011,32'b0111110110011001110011110000100,32'b0111110100100101111010011101001,32'b0111101100101101110001111001010,32'b0111111000000000110000101101101,32'b1111111000111010000010000001010,32'b1111101101010101111100011101101,32'b1111101000111111010001001111001,32'b1111110100111110101110011111111,32'b0111110110111100011100111100100,32'b0111111001101010010111010111000,32'b0111111010100101100001011100110,32'b1111100101000001110101011000101,32'b0111111000001011100110010010101,32'b0111011110110001111101100010000,32'b0111111001111100001110001100101,32'b1111110101101010101011010101101,32'b1111111001111110011011111000000,32'b1111101001000010110100001011111,32'b0111110101110100011010100001100,32'b0111111010110111111110000111011,32'b0111111010011000101100011110101,32'b1111111000101000011010001111110,32'b0111111011101001010110001111010,32'b1111110110010101110101001101100,32'b1111111011000001100101010000110,32'b1111101011100000001000000010101,32'b0111111000011100011100010010001,32'b1111111001110000011000110110000,32'b1111111001001110101100000010010,32'b1111110001100100110010111000110,32'b1111110101110011011100010000000,32'b0111110100111110001110011100011,32'b0111111010100111111110101100000,32'b0111111001100011110111111100100,32'b0111111010110000110100000111010,32'b0111110101011100110001100101010,32'b1111110111101111111010010011001,32'b1111110100100011001001010111010,32'b1111111011110010110001010101100,32'b1111110010101110011000111110111,32'b0111110011101011101001001000101,32'b0111111010001111111001011011101,32'b1111110100010100011111111100011,32'b1111111001011101111110010010101,32'b1111110100000010111000011101000,32'b1111110011011110010110101010010,32'b0111110100100010100100001101000,32'b1111110110011100100011011001100,32'b0111110111111100100010010011010,32'b0111111000001001110101010011011,32'b1111110010101101110100010111110,32'b0111101011111101111000111111110,32'b1111111000010101111110111101001,32'b0111111010011111011100001000011,32'b0111110101110100011000100111000,32'b0111110011001100001010000111010,32'b1111111001100000001100100101001,32'b1111110101010000001000100011101,32'b1111100010110111010110101010100,32'b0111110001001101100110001110000,32'b1111110011111000000010010000100,32'b0111111010110111010111100011010,32'b0111101110011110110110001011110,32'b0111110001011011000101010010011,32'b1111111001001110101001101111110,32'b0111110101010101111001000000000,32'b0111111011011101011011000100111,32'b0111110101000111000101000000101,32'b1111110000000111111000101000001,32'b0111100101000100111010101000110,32'b0111111011111100101000101100100,32'b1111111011010111011010101101100,32'b1111111000100010111110110111110,32'b0111110101101111010100011000111};
    assign bias = {32'b1111101011101010001110010000110,32'b1110111101111000000101010000000,32'b0111101011010011001100101101011,32'b1111011110000110010001011000000,32'b1111010111100010100011111100001,32'b0111100101000101001001011010100,32'b1111001111000000110010100111110,32'b1111101000110000000001010110010};
endmodule